`timescale 1ns / 1ps
/* --------------------------------- */
/* YOUR DUT IMPLEMENTATION GOES HERE */
/* --------------------------------- */

// module dut_test #(
//     parameter IN_BUS_WIDTH = 256,
//     parameter OUT_BUS_WIDTH = 256
// )(
//     input logic     clk,
//     input logic     rst_n,
//     input logic     [IN_BUS_WIDTH-1:0] in,
//     output logic    [OUT_BUS_WIDTH-1:0] out
// );

// ...
    
// endmodule
